library verilog;
use verilog.vl_types.all;
entity tb_n is
end tb_n;
