-- megafunction wizard: %LPM_MULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mult 

-- ============================================================
-- File Name: altera_mult_30b.vhd
-- Megafunction Name(s):
-- 			lpm_mult
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.all;

ENTITY altera_mult_30b IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (29 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (29 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (60 DOWNTO 0)
	);
END altera_mult_30b;


ARCHITECTURE SYN OF altera_mult_30b IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (60 DOWNTO 0);



	COMPONENT lpm_mult
	GENERIC (
		lpm_hint		: STRING;
		lpm_pipeline		: NATURAL;
		lpm_representation		: STRING;
		lpm_type		: STRING;
		lpm_widtha		: NATURAL;
		lpm_widthb		: NATURAL;
		lpm_widthp		: NATURAL
	);
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (29 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (29 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (60 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(60 DOWNTO 0);

	lpm_mult_component : lpm_mult
	GENERIC MAP (
		lpm_hint => "MAXIMIZE_SPEED=5",
		lpm_pipeline => 1,
		lpm_representation => "SIGNED",
		lpm_type => "LPM_MULT",
		lpm_widtha => 30,
		lpm_widthb => 30,
		lpm_widthp => 61
	)
	PORT MAP (
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: AutoSizeResult NUMERIC "0"
-- Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
-- Retrieval info: PRIVATE: ConstantB NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "1"
-- Retrieval info: PRIVATE: Latency NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: SignedMult NUMERIC "1"
-- Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
-- Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
-- Retrieval info: PRIVATE: WidthA NUMERIC "30"
-- Retrieval info: PRIVATE: WidthB NUMERIC "30"
-- Retrieval info: PRIVATE: WidthP NUMERIC "61"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: PRIVATE: optimize NUMERIC "0"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=5"
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
-- Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "30"
-- Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "30"
-- Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "61"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 30 0 INPUT NODEFVAL "dataa[29..0]"
-- Retrieval info: USED_PORT: datab 0 0 30 0 INPUT NODEFVAL "datab[29..0]"
-- Retrieval info: USED_PORT: result 0 0 61 0 OUTPUT NODEFVAL "result[60..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 30 0 dataa 0 0 30 0
-- Retrieval info: CONNECT: @datab 0 0 30 0 datab 0 0 30 0
-- Retrieval info: CONNECT: result 0 0 61 0 @result 0 0 61 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altera_mult_30b.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altera_mult_30b.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altera_mult_30b.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altera_mult_30b.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altera_mult_30b_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
