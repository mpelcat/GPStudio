/* Dual-core ARM Cortex-A9 instance (wrapper for Qsys generation) */
module arm
(
		input  wire        clk_proc,                           
		input  wire        reset_reset_n,                         
		output wire [14:0] memory_mem_a,                          
		output wire [2:0]  memory_mem_ba,                         
		output wire        memory_mem_ck,                         
		output wire        memory_mem_ck_n,                       
		output wire        memory_mem_cke,                        
		output wire        memory_mem_cs_n,                       
		output wire        memory_mem_ras_n,                      
		output wire        memory_mem_cas_n,                      
		output wire        memory_mem_we_n,                       
		output wire        memory_mem_reset_n,                    
		inout  wire [31:0] memory_mem_dq,                         
		inout  wire [3:0]  memory_mem_dqs,                        
		inout  wire [3:0]  memory_mem_dqs_n,                      
		output wire        memory_mem_odt,                        
		output wire [3:0]  memory_mem_dm,                         
		input  wire        memory_oct_rzqin,                      
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, 
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, 
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, 
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, 
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,     
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,     
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,     
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,     
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,     
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,     
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     
		output wire        hps_0_hps_io_hps_io_spim0_inst_CLK,    
		output wire        hps_0_hps_io_hps_io_spim0_inst_MOSI,   
		input  wire        hps_0_hps_io_hps_io_spim0_inst_MISO,   
		output wire        hps_0_hps_io_hps_io_spim0_inst_SS0,    
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,    
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,   
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,   
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,    
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,     
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,     
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO00,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO55,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO56,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO62,  
		output wire        hps_0_h2f_reset_reset_n,               
		input  wire        hps_0_f2h_cold_reset_req_reset_n,      
		input  wire        hps_0_f2h_debug_reset_req_reset_n,     
		input  wire        hps_0_f2h_warm_reset_req_reset_n,      
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,  
		output wire        out0_fv,                               
		output wire        out0_dv,                               
		output wire [OUT0_SIZE-1:0] out0_data,                             
		output wire        out1_fv,                               
		output wire        out1_dv,                               
		output wire [OUT1_SIZE-1:0] out1_data,                             
		input  wire        in0_dv,                                
		input  wire [IN0_SIZE-1:0] in0_data,                              
		input  wire        in0_fv,                                
		input  wire        in1_dv,                                
		input  wire [IN1_SIZE-1:0] in1_data,                              
		input  wire        in1_fv,                                
		output wire [MASTER_ADDR_WIDTH-1:0]  master_addr_o,                         
		output wire        master_wr_o,                           
		output wire        master_rd_o,                           
		output wire [31:0] master_datawr_o,                       
		input  wire [31:0] master_datard_i,                       
		input  wire        master_waitreq

);

parameter CLK_PROC_FREQ = 50000000;
parameter CLK_CLK_FREQ 	= 50000000;
parameter IN0_SIZE		= 16;
parameter IN1_SIZE		= 16;
parameter OUT0_SIZE		= 16;
parameter OUT1_SIZE		= 16;
parameter MASTER_ADDR_WIDTH = 32;

soc_system soc_system_inst
(
		.clk_clk(clk_proc),
		.reset_reset_n(reset_reset_n),
		.memory_mem_a(memory_mem_a),
		.memory_mem_ba(memory_mem_ba),
		.memory_mem_ck(memory_mem_ck),
		.memory_mem_ck_n(memory_mem_ck_n),
		.memory_mem_cke(memory_mem_cke),
		.memory_mem_cs_n(memory_mem_cs_n),
		.memory_mem_ras_n(memory_mem_ras_n),
		.memory_mem_cas_n(memory_mem_cas_n),
		.memory_mem_we_n(memory_mem_we_n),
		.memory_mem_reset_n(memory_mem_reset_n),
		.memory_mem_dq(memory_mem_dq),
		.memory_mem_dqs(memory_mem_dqs),
		.memory_mem_dqs_n(memory_mem_dqs_n),
		.memory_mem_odt(memory_mem_odt),
		.memory_mem_dm(memory_mem_dm),
		.memory_oct_rzqin(memory_oct_rzqin),
		.hps_0_hps_io_hps_io_emac1_inst_TX_CLK(hps_0_hps_io_hps_io_emac1_inst_TX_CLK),
		.hps_0_hps_io_hps_io_emac1_inst_TXD0(hps_0_hps_io_hps_io_emac1_inst_TXD0),
		.hps_0_hps_io_hps_io_emac1_inst_TXD1(hps_0_hps_io_hps_io_emac1_inst_TXD1),
		.hps_0_hps_io_hps_io_emac1_inst_TXD2(hps_0_hps_io_hps_io_emac1_inst_TXD2),
		.hps_0_hps_io_hps_io_emac1_inst_TXD3(hps_0_hps_io_hps_io_emac1_inst_TXD3),
		.hps_0_hps_io_hps_io_emac1_inst_RXD0(hps_0_hps_io_hps_io_emac1_inst_RXD0),
		.hps_0_hps_io_hps_io_emac1_inst_MDIO(hps_0_hps_io_hps_io_emac1_inst_MDIO),
		.hps_0_hps_io_hps_io_emac1_inst_MDC(hps_0_hps_io_hps_io_emac1_inst_MDC),
		.hps_0_hps_io_hps_io_emac1_inst_RX_CTL(hps_0_hps_io_hps_io_emac1_inst_RX_CTL),
		.hps_0_hps_io_hps_io_emac1_inst_TX_CTL(hps_0_hps_io_hps_io_emac1_inst_TX_CTL),
		.hps_0_hps_io_hps_io_emac1_inst_RX_CLK(hps_0_hps_io_hps_io_emac1_inst_RX_CLK),
		.hps_0_hps_io_hps_io_emac1_inst_RXD1(hps_0_hps_io_hps_io_emac1_inst_RXD1),
		.hps_0_hps_io_hps_io_emac1_inst_RXD2(hps_0_hps_io_hps_io_emac1_inst_RXD2),
		.hps_0_hps_io_hps_io_emac1_inst_RXD3(hps_0_hps_io_hps_io_emac1_inst_RXD3),
		.hps_0_hps_io_hps_io_qspi_inst_IO0(hps_0_hps_io_hps_io_qspi_inst_IO0),
		.hps_0_hps_io_hps_io_qspi_inst_IO1(hps_0_hps_io_hps_io_qspi_inst_IO1),
		.hps_0_hps_io_hps_io_qspi_inst_IO2(hps_0_hps_io_hps_io_qspi_inst_IO2),
		.hps_0_hps_io_hps_io_qspi_inst_IO3(hps_0_hps_io_hps_io_qspi_inst_IO3),
		.hps_0_hps_io_hps_io_qspi_inst_SS0(hps_0_hps_io_hps_io_qspi_inst_SS0),
		.hps_0_hps_io_hps_io_qspi_inst_CLK(hps_0_hps_io_hps_io_qspi_inst_CLK),
		.hps_0_hps_io_hps_io_sdio_inst_CMD(hps_0_hps_io_hps_io_sdio_inst_CMD),
		.hps_0_hps_io_hps_io_sdio_inst_D0(hps_0_hps_io_hps_io_sdio_inst_D0),
		.hps_0_hps_io_hps_io_sdio_inst_D1(hps_0_hps_io_hps_io_sdio_inst_D1),
		.hps_0_hps_io_hps_io_sdio_inst_CLK(hps_0_hps_io_hps_io_sdio_inst_CLK),
		.hps_0_hps_io_hps_io_sdio_inst_D2(hps_0_hps_io_hps_io_sdio_inst_D2),
		.hps_0_hps_io_hps_io_sdio_inst_D3(hps_0_hps_io_hps_io_sdio_inst_D3),
		.hps_0_hps_io_hps_io_usb1_inst_D0(hps_0_hps_io_hps_io_usb1_inst_D0),
		.hps_0_hps_io_hps_io_usb1_inst_D1(hps_0_hps_io_hps_io_usb1_inst_D1),
		.hps_0_hps_io_hps_io_usb1_inst_D2(hps_0_hps_io_hps_io_usb1_inst_D2),
		.hps_0_hps_io_hps_io_usb1_inst_D3(hps_0_hps_io_hps_io_usb1_inst_D3),
		.hps_0_hps_io_hps_io_usb1_inst_D4(hps_0_hps_io_hps_io_usb1_inst_D4),
		.hps_0_hps_io_hps_io_usb1_inst_D5(hps_0_hps_io_hps_io_usb1_inst_D5),
		.hps_0_hps_io_hps_io_usb1_inst_D6(hps_0_hps_io_hps_io_usb1_inst_D6),
		.hps_0_hps_io_hps_io_usb1_inst_D7(hps_0_hps_io_hps_io_usb1_inst_D7),
		.hps_0_hps_io_hps_io_usb1_inst_CLK(hps_0_hps_io_hps_io_usb1_inst_CLK),
		.hps_0_hps_io_hps_io_usb1_inst_STP(hps_0_hps_io_hps_io_usb1_inst_STP),
		.hps_0_hps_io_hps_io_usb1_inst_DIR(hps_0_hps_io_hps_io_usb1_inst_DIR),
		.hps_0_hps_io_hps_io_usb1_inst_NXT(hps_0_hps_io_hps_io_usb1_inst_NXT),
		.hps_0_hps_io_hps_io_spim0_inst_CLK(hps_0_hps_io_hps_io_spim0_inst_CLK),
		.hps_0_hps_io_hps_io_spim0_inst_MOSI(hps_0_hps_io_hps_io_spim0_inst_MOSI),
		.hps_0_hps_io_hps_io_spim0_inst_MISO(hps_0_hps_io_hps_io_spim0_inst_MISO),
		.hps_0_hps_io_hps_io_spim0_inst_SS0(hps_0_hps_io_hps_io_spim0_inst_SS0),
		.hps_0_hps_io_hps_io_spim1_inst_CLK(hps_0_hps_io_hps_io_spim1_inst_CLK),
		.hps_0_hps_io_hps_io_spim1_inst_MOSI(hps_0_hps_io_hps_io_spim1_inst_MOSI),
		.hps_0_hps_io_hps_io_spim1_inst_MISO(hps_0_hps_io_hps_io_spim1_inst_MISO),
		.hps_0_hps_io_hps_io_spim1_inst_SS0(hps_0_hps_io_hps_io_spim1_inst_SS0),
		.hps_0_hps_io_hps_io_uart0_inst_RX(hps_0_hps_io_hps_io_uart0_inst_RX),
		.hps_0_hps_io_hps_io_uart0_inst_TX(hps_0_hps_io_hps_io_uart0_inst_TX),
		.hps_0_hps_io_hps_io_i2c1_inst_SDA(hps_0_hps_io_hps_io_i2c1_inst_SDA),
		.hps_0_hps_io_hps_io_i2c1_inst_SCL(hps_0_hps_io_hps_io_i2c1_inst_SCL),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO00(hps_0_hps_io_hps_io_gpio_inst_GPIO00),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO09(hps_0_hps_io_hps_io_gpio_inst_GPIO09),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO35(hps_0_hps_io_hps_io_gpio_inst_GPIO35),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO48(hps_0_hps_io_hps_io_gpio_inst_GPIO48),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO53(hps_0_hps_io_hps_io_gpio_inst_GPIO53),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO54(hps_0_hps_io_hps_io_gpio_inst_GPIO54),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO55(hps_0_hps_io_hps_io_gpio_inst_GPIO55),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO56(hps_0_hps_io_hps_io_gpio_inst_GPIO56),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO61(hps_0_hps_io_hps_io_gpio_inst_GPIO61),
		.hps_0_hps_io_hps_io_gpio_inst_GPIO62(hps_0_hps_io_hps_io_gpio_inst_GPIO62),
		.hps_0_h2f_reset_reset_n(hps_0_h2f_reset_reset_n),
		.hps_0_f2h_cold_reset_req_reset_n(hps_0_f2h_cold_reset_req_reset_n),
		.hps_0_f2h_debug_reset_req_reset_n(hps_0_f2h_debug_reset_req_reset_n),
		.hps_0_f2h_warm_reset_req_reset_n(hps_0_f2h_warm_reset_req_reset_n),
		.hps_0_f2h_stm_hw_events_stm_hwevents(hps_0_f2h_stm_hw_events_stm_hwevents),
		.out0_fv(out0_fv),
		.out0_dv(out0_dv),
		.out0_data(out0_data),
		.out1_fv(out1_fv),
		.out1_dv(out1_dv),
		.out1_data(out1_data),
		.in0_dv(in0_dv),
		.in0_data(in0_data),
		.in0_fv(in0_fv),
		.in1_dv(in1_dv),
		.in1_data(in1_data),
		.in1_fv(in1_fv),
		.master_addr_o(master_addr_o),
		.master_wr_o(master_wr_o),
		.master_rd_o(master_rd_o),
		.master_datawr_o(master_datawr_o),
		.master_datard_i(master_datard_i),
		.master_waitreq(master_waitreq)
);

endmodule
